package TestbenchClasses;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "AxisWord.sv"
    `include "MasterMonitor.sv"
    `include "MasterDriver.sv"
    `include "RandomPacket.sv"
    `include "MasterAgent.sv"
    `include "PacketSequence.sv"
    `include "SlaveMonitor.sv"
    `include "SlaveDriver.sv"
    `include "SlaveAgent.sv"
    `include "Scoreboard.sv"
    `include "Environment.sv"
    `include "random_test.sv"
endpackage
